module grass_sprite(
    input wire clk,
    input wire [4:0] pixel_x,      
    input wire [4:0] pixel_y,      
    output reg [5:0] pixel_color   
);

    reg [8:0] sprite_memory [0:1023];  

    wire [9:0] pixel_index = {pixel_y, pixel_x}; 

    initial begin
        sprite_memory[0] = 6'b00_00_00;
        sprite_memory[1] = 6'b00_00_00;
        sprite_memory[2] = 6'b11_01_00;
        sprite_memory[3] = 6'b11_01_00;
        sprite_memory[4] = 6'b11_01_00;
        sprite_memory[5] = 6'b11_01_00;
        sprite_memory[6] = 6'b11_01_00;
        sprite_memory[7] = 6'b11_01_00;
        sprite_memory[8] = 6'b11_01_00;
        sprite_memory[9] = 6'b11_01_00;
        sprite_memory[10] = 6'b11_01_00;
        sprite_memory[11] = 6'b11_01_00;
        sprite_memory[12] = 6'b11_01_00;
        sprite_memory[13] = 6'b11_01_00;
        sprite_memory[14] = 6'b11_01_00;
        sprite_memory[15] = 6'b11_01_00;
        sprite_memory[16] = 6'b11_01_00;
        sprite_memory[17] = 6'b11_01_00;
        sprite_memory[18] = 6'b11_01_00;
        sprite_memory[19] = 6'b11_01_00;
        sprite_memory[20] = 6'b11_01_00;
        sprite_memory[21] = 6'b11_01_00;
        sprite_memory[22] = 6'b11_01_00;
        sprite_memory[23] = 6'b11_01_00;
        sprite_memory[24] = 6'b11_01_00;
        sprite_memory[25] = 6'b11_01_00;
        sprite_memory[26] = 6'b11_01_00;
        sprite_memory[27] = 6'b11_01_00;
        sprite_memory[28] = 6'b11_01_00;
        sprite_memory[29] = 6'b11_01_00;
        sprite_memory[30] = 6'b11_01_00;
        sprite_memory[31] = 6'b11_01_00;
        sprite_memory[32] = 6'b00_00_00;
        sprite_memory[33] = 6'b00_00_00;
        sprite_memory[34] = 6'b11_01_00;
        sprite_memory[35] = 6'b11_01_00;
        sprite_memory[36] = 6'b11_01_00;
        sprite_memory[37] = 6'b11_01_00;
        sprite_memory[38] = 6'b11_01_00;
        sprite_memory[39] = 6'b11_01_00;
        sprite_memory[40] = 6'b11_01_00;
        sprite_memory[41] = 6'b11_01_00;
        sprite_memory[42] = 6'b11_01_00;
        sprite_memory[43] = 6'b11_01_00;
        sprite_memory[44] = 6'b11_01_00;
        sprite_memory[45] = 6'b00_00_00;
        sprite_memory[46] = 6'b11_01_00;
        sprite_memory[47] = 6'b11_01_00;
        sprite_memory[48] = 6'b11_01_00;
        sprite_memory[49] = 6'b11_01_00;
        sprite_memory[50] = 6'b11_01_00;
        sprite_memory[51] = 6'b11_01_00;
        sprite_memory[52] = 6'b11_01_00;
        sprite_memory[53] = 6'b11_01_00;
        sprite_memory[54] = 6'b11_01_00;
        sprite_memory[55] = 6'b11_01_00;
        sprite_memory[56] = 6'b11_01_00;
        sprite_memory[57] = 6'b11_01_00;
        sprite_memory[58] = 6'b11_01_00;
        sprite_memory[59] = 6'b11_01_00;
        sprite_memory[60] = 6'b11_01_00;
        sprite_memory[61] = 6'b11_01_00;
        sprite_memory[62] = 6'b11_01_00;
        sprite_memory[63] = 6'b11_01_00;
        sprite_memory[64] = 6'b00_00_00;
        sprite_memory[65] = 6'b11_01_00;
        sprite_memory[66] = 6'b11_01_00;
        sprite_memory[67] = 6'b11_01_00;
        sprite_memory[68] = 6'b11_01_00;
        sprite_memory[69] = 6'b11_01_00;
        sprite_memory[70] = 6'b00_00_00;
        sprite_memory[71] = 6'b11_01_00;
        sprite_memory[72] = 6'b11_01_00;
        sprite_memory[73] = 6'b11_01_00;
        sprite_memory[74] = 6'b11_01_00;
        sprite_memory[75] = 6'b11_01_00;
        sprite_memory[76] = 6'b11_01_00;
        sprite_memory[77] = 6'b10_01_01;
        sprite_memory[78] = 6'b00_00_00;
        sprite_memory[79] = 6'b11_01_00;
        sprite_memory[80] = 6'b11_01_00;
        sprite_memory[81] = 6'b11_01_00;
        sprite_memory[82] = 6'b11_01_00;
        sprite_memory[83] = 6'b11_01_00;
        sprite_memory[84] = 6'b11_01_00;
        sprite_memory[85] = 6'b11_01_00;
        sprite_memory[86] = 6'b11_01_00;
        sprite_memory[87] = 6'b11_01_00;
        sprite_memory[88] = 6'b11_01_00;
        sprite_memory[89] = 6'b11_01_00;
        sprite_memory[90] = 6'b11_01_00;
        sprite_memory[91] = 6'b00_00_00;
        sprite_memory[92] = 6'b11_01_00;
        sprite_memory[93] = 6'b11_01_00;
        sprite_memory[94] = 6'b11_01_00;
        sprite_memory[95] = 6'b11_01_00;
        sprite_memory[96] = 6'b00_00_00;
        sprite_memory[97] = 6'b11_01_00;
        sprite_memory[98] = 6'b11_01_00;
        sprite_memory[99] = 6'b11_01_00;
        sprite_memory[100] = 6'b11_01_00;
        sprite_memory[101] = 6'b11_01_00;
        sprite_memory[102] = 6'b11_01_00;
        sprite_memory[103] = 6'b11_01_00;
        sprite_memory[104] = 6'b11_01_00;
        sprite_memory[105] = 6'b11_01_00;
        sprite_memory[106] = 6'b11_01_00;
        sprite_memory[107] = 6'b11_01_00;
        sprite_memory[108] = 6'b11_01_00;
        sprite_memory[109] = 6'b10_01_01;
        sprite_memory[110] = 6'b11_01_00;
        sprite_memory[111] = 6'b11_01_00;
        sprite_memory[112] = 6'b11_01_00;
        sprite_memory[113] = 6'b11_01_00;
        sprite_memory[114] = 6'b11_01_00;
        sprite_memory[115] = 6'b11_01_00;
        sprite_memory[116] = 6'b11_01_00;
        sprite_memory[117] = 6'b11_01_00;
        sprite_memory[118] = 6'b00_00_00;
        sprite_memory[119] = 6'b11_01_00;
        sprite_memory[120] = 6'b11_01_00;
        sprite_memory[121] = 6'b11_01_00;
        sprite_memory[122] = 6'b11_01_00;
        sprite_memory[123] = 6'b10_01_01;
        sprite_memory[124] = 6'b00_00_00;
        sprite_memory[125] = 6'b11_01_00;
        sprite_memory[126] = 6'b11_01_00;
        sprite_memory[127] = 6'b11_01_00;
        sprite_memory[128] = 6'b00_00_00;
        sprite_memory[129] = 6'b11_01_00;
        sprite_memory[130] = 6'b11_01_00;
        sprite_memory[131] = 6'b00_00_00;
        sprite_memory[132] = 6'b11_01_00;
        sprite_memory[133] = 6'b11_01_00;
        sprite_memory[134] = 6'b11_01_00;
        sprite_memory[135] = 6'b11_01_00;
        sprite_memory[136] = 6'b11_01_00;
        sprite_memory[137] = 6'b11_01_00;
        sprite_memory[138] = 6'b11_01_00;
        sprite_memory[139] = 6'b11_01_00;
        sprite_memory[140] = 6'b11_01_00;
        sprite_memory[141] = 6'b11_01_00;
        sprite_memory[142] = 6'b11_01_00;
        sprite_memory[143] = 6'b11_01_00;
        sprite_memory[144] = 6'b11_01_00;
        sprite_memory[145] = 6'b11_01_00;
        sprite_memory[146] = 6'b11_01_00;
        sprite_memory[147] = 6'b11_01_00;
        sprite_memory[148] = 6'b11_01_00;
        sprite_memory[149] = 6'b11_01_00;
        sprite_memory[150] = 6'b11_01_00;
        sprite_memory[151] = 6'b11_01_00;
        sprite_memory[152] = 6'b11_01_00;
        sprite_memory[153] = 6'b11_01_00;
        sprite_memory[154] = 6'b11_01_00;
        sprite_memory[155] = 6'b10_01_01;
        sprite_memory[156] = 6'b11_01_00;
        sprite_memory[157] = 6'b11_01_00;
        sprite_memory[158] = 6'b11_01_00;
        sprite_memory[159] = 6'b11_01_00;
        sprite_memory[160] = 6'b00_00_00;
        sprite_memory[161] = 6'b11_01_00;
        sprite_memory[162] = 6'b11_01_00;
        sprite_memory[163] = 6'b10_01_01;
        sprite_memory[164] = 6'b00_00_00;
        sprite_memory[165] = 6'b11_01_00;
        sprite_memory[166] = 6'b11_01_00;
        sprite_memory[167] = 6'b11_01_00;
        sprite_memory[168] = 6'b11_01_00;
        sprite_memory[169] = 6'b11_01_00;
        sprite_memory[170] = 6'b11_01_00;
        sprite_memory[171] = 6'b11_01_00;
        sprite_memory[172] = 6'b11_01_00;
        sprite_memory[173] = 6'b11_01_00;
        sprite_memory[174] = 6'b11_01_00;
        sprite_memory[175] = 6'b00_00_00;
        sprite_memory[176] = 6'b11_01_00;
        sprite_memory[177] = 6'b11_01_00;
        sprite_memory[178] = 6'b11_01_00;
        sprite_memory[179] = 6'b11_01_00;
        sprite_memory[180] = 6'b00_00_00;
        sprite_memory[181] = 6'b11_01_00;
        sprite_memory[182] = 6'b11_01_00;
        sprite_memory[183] = 6'b11_01_00;
        sprite_memory[184] = 6'b11_01_00;
        sprite_memory[185] = 6'b11_01_00;
        sprite_memory[186] = 6'b11_01_00;
        sprite_memory[187] = 6'b11_01_00;
        sprite_memory[188] = 6'b11_01_00;
        sprite_memory[189] = 6'b11_01_00;
        sprite_memory[190] = 6'b11_01_00;
        sprite_memory[191] = 6'b11_01_00;
        sprite_memory[192] = 6'b00_00_00;
        sprite_memory[193] = 6'b11_01_00;
        sprite_memory[194] = 6'b11_01_00;
        sprite_memory[195] = 6'b10_01_01;
        sprite_memory[196] = 6'b11_01_00;
        sprite_memory[197] = 6'b11_01_00;
        sprite_memory[198] = 6'b11_01_00;
        sprite_memory[199] = 6'b11_01_00;
        sprite_memory[200] = 6'b11_01_00;
        sprite_memory[201] = 6'b00_00_00;
        sprite_memory[202] = 6'b11_01_00;
        sprite_memory[203] = 6'b11_01_00;
        sprite_memory[204] = 6'b11_01_00;
        sprite_memory[205] = 6'b11_01_00;
        sprite_memory[206] = 6'b11_01_00;
        sprite_memory[207] = 6'b11_01_00;
        sprite_memory[208] = 6'b11_01_00;
        sprite_memory[209] = 6'b11_01_00;
        sprite_memory[210] = 6'b11_01_00;
        sprite_memory[211] = 6'b11_01_00;
        sprite_memory[212] = 6'b10_01_01;
        sprite_memory[213] = 6'b00_00_00;
        sprite_memory[214] = 6'b11_01_00;
        sprite_memory[215] = 6'b11_01_00;
        sprite_memory[216] = 6'b11_01_00;
        sprite_memory[217] = 6'b11_01_00;
        sprite_memory[218] = 6'b11_01_00;
        sprite_memory[219] = 6'b11_01_00;
        sprite_memory[220] = 6'b11_01_00;
        sprite_memory[221] = 6'b11_01_00;
        sprite_memory[222] = 6'b11_01_00;
        sprite_memory[223] = 6'b11_01_00;
        sprite_memory[224] = 6'b00_00_00;
        sprite_memory[225] = 6'b00_00_00;
        sprite_memory[226] = 6'b11_01_00;
        sprite_memory[227] = 6'b11_01_00;
        sprite_memory[228] = 6'b11_01_00;
        sprite_memory[229] = 6'b11_01_00;
        sprite_memory[230] = 6'b11_01_00;
        sprite_memory[231] = 6'b11_01_00;
        sprite_memory[232] = 6'b11_01_00;
        sprite_memory[233] = 6'b10_01_01;
        sprite_memory[234] = 6'b00_00_00;
        sprite_memory[235] = 6'b11_01_00;
        sprite_memory[236] = 6'b11_01_00;
        sprite_memory[237] = 6'b11_01_00;
        sprite_memory[238] = 6'b11_01_00;
        sprite_memory[239] = 6'b11_01_00;
        sprite_memory[240] = 6'b11_01_00;
        sprite_memory[241] = 6'b11_01_00;
        sprite_memory[242] = 6'b11_01_00;
        sprite_memory[243] = 6'b11_01_00;
        sprite_memory[244] = 6'b10_01_01;
        sprite_memory[245] = 6'b11_01_00;
        sprite_memory[246] = 6'b11_01_00;
        sprite_memory[247] = 6'b11_01_00;
        sprite_memory[248] = 6'b11_01_00;
        sprite_memory[249] = 6'b11_01_00;
        sprite_memory[250] = 6'b11_01_00;
        sprite_memory[251] = 6'b11_01_00;
        sprite_memory[252] = 6'b00_00_00;
        sprite_memory[253] = 6'b11_01_00;
        sprite_memory[254] = 6'b11_01_00;
        sprite_memory[255] = 6'b11_01_00;
        sprite_memory[256] = 6'b00_00_00;
        sprite_memory[257] = 6'b00_00_00;
        sprite_memory[258] = 6'b00_00_00;
        sprite_memory[259] = 6'b11_01_00;
        sprite_memory[260] = 6'b11_01_00;
        sprite_memory[261] = 6'b11_01_00;
        sprite_memory[262] = 6'b11_01_00;
        sprite_memory[263] = 6'b11_01_00;
        sprite_memory[264] = 6'b11_01_00;
        sprite_memory[265] = 6'b10_01_01;
        sprite_memory[266] = 6'b11_01_00;
        sprite_memory[267] = 6'b11_01_00;
        sprite_memory[268] = 6'b11_01_00;
        sprite_memory[269] = 6'b11_01_00;
        sprite_memory[270] = 6'b11_01_00;
        sprite_memory[271] = 6'b11_01_00;
        sprite_memory[272] = 6'b11_01_00;
        sprite_memory[273] = 6'b11_01_00;
        sprite_memory[274] = 6'b11_01_00;
        sprite_memory[275] = 6'b11_01_00;
        sprite_memory[276] = 6'b11_01_00;
        sprite_memory[277] = 6'b11_01_00;
        sprite_memory[278] = 6'b11_01_00;
        sprite_memory[279] = 6'b11_01_00;
        sprite_memory[280] = 6'b11_01_00;
        sprite_memory[281] = 6'b11_01_00;
        sprite_memory[282] = 6'b11_01_00;
        sprite_memory[283] = 6'b11_01_00;
        sprite_memory[284] = 6'b10_01_01;
        sprite_memory[285] = 6'b00_00_00;
        sprite_memory[286] = 6'b11_01_00;
        sprite_memory[287] = 6'b11_01_00;
        sprite_memory[288] = 6'b00_00_00;
        sprite_memory[289] = 6'b00_00_00;
        sprite_memory[290] = 6'b11_01_00;
        sprite_memory[291] = 6'b11_01_00;
        sprite_memory[292] = 6'b11_01_00;
        sprite_memory[293] = 6'b11_01_00;
        sprite_memory[294] = 6'b11_01_00;
        sprite_memory[295] = 6'b11_01_00;
        sprite_memory[296] = 6'b11_01_00;
        sprite_memory[297] = 6'b11_01_00;
        sprite_memory[298] = 6'b11_01_00;
        sprite_memory[299] = 6'b11_01_00;
        sprite_memory[300] = 6'b11_01_00;
        sprite_memory[301] = 6'b11_01_00;
        sprite_memory[302] = 6'b11_01_00;
        sprite_memory[303] = 6'b11_01_00;
        sprite_memory[304] = 6'b00_00_00;
        sprite_memory[305] = 6'b11_01_00;
        sprite_memory[306] = 6'b11_01_00;
        sprite_memory[307] = 6'b11_01_00;
        sprite_memory[308] = 6'b11_01_00;
        sprite_memory[309] = 6'b11_01_00;
        sprite_memory[310] = 6'b11_01_00;
        sprite_memory[311] = 6'b11_01_00;
        sprite_memory[312] = 6'b11_01_00;
        sprite_memory[313] = 6'b11_01_00;
        sprite_memory[314] = 6'b11_01_00;
        sprite_memory[315] = 6'b11_01_00;
        sprite_memory[316] = 6'b10_01_01;
        sprite_memory[317] = 6'b11_01_00;
        sprite_memory[318] = 6'b11_01_00;
        sprite_memory[319] = 6'b00_00_00;
        sprite_memory[320] = 6'b00_00_00;
        sprite_memory[321] = 6'b11_01_00;
        sprite_memory[322] = 6'b11_01_00;
        sprite_memory[323] = 6'b11_01_00;
        sprite_memory[324] = 6'b11_01_00;
        sprite_memory[325] = 6'b11_01_00;
        sprite_memory[326] = 6'b11_01_00;
        sprite_memory[327] = 6'b11_01_00;
        sprite_memory[328] = 6'b11_01_00;
        sprite_memory[329] = 6'b11_01_00;
        sprite_memory[330] = 6'b11_01_00;
        sprite_memory[331] = 6'b11_01_00;
        sprite_memory[332] = 6'b11_01_00;
        sprite_memory[333] = 6'b11_01_00;
        sprite_memory[334] = 6'b11_01_00;
        sprite_memory[335] = 6'b11_01_00;
        sprite_memory[336] = 6'b10_01_01;
        sprite_memory[337] = 6'b00_00_00;
        sprite_memory[338] = 6'b11_01_00;
        sprite_memory[339] = 6'b11_01_00;
        sprite_memory[340] = 6'b11_01_00;
        sprite_memory[341] = 6'b11_01_00;
        sprite_memory[342] = 6'b11_01_00;
        sprite_memory[343] = 6'b11_01_00;
        sprite_memory[344] = 6'b11_01_00;
        sprite_memory[345] = 6'b00_00_00;
        sprite_memory[346] = 6'b11_01_00;
        sprite_memory[347] = 6'b11_01_00;
        sprite_memory[348] = 6'b11_01_00;
        sprite_memory[349] = 6'b11_01_00;
        sprite_memory[350] = 6'b11_01_00;
        sprite_memory[351] = 6'b00_00_00;
        sprite_memory[352] = 6'b00_00_00;
        sprite_memory[353] = 6'b11_01_00;
        sprite_memory[354] = 6'b11_01_00;
        sprite_memory[355] = 6'b11_01_00;
        sprite_memory[356] = 6'b11_01_00;
        sprite_memory[357] = 6'b11_01_00;
        sprite_memory[358] = 6'b11_01_00;
        sprite_memory[359] = 6'b11_01_00;
        sprite_memory[360] = 6'b11_01_00;
        sprite_memory[361] = 6'b11_01_00;
        sprite_memory[362] = 6'b11_01_00;
        sprite_memory[363] = 6'b11_01_00;
        sprite_memory[364] = 6'b11_01_00;
        sprite_memory[365] = 6'b11_01_00;
        sprite_memory[366] = 6'b11_01_00;
        sprite_memory[367] = 6'b11_01_00;
        sprite_memory[368] = 6'b10_01_01;
        sprite_memory[369] = 6'b11_01_00;
        sprite_memory[370] = 6'b11_01_00;
        sprite_memory[371] = 6'b11_01_00;
        sprite_memory[372] = 6'b11_01_00;
        sprite_memory[373] = 6'b11_01_00;
        sprite_memory[374] = 6'b11_01_00;
        sprite_memory[375] = 6'b11_01_00;
        sprite_memory[376] = 6'b11_01_00;
        sprite_memory[377] = 6'b11_01_00;
        sprite_memory[378] = 6'b11_01_00;
        sprite_memory[379] = 6'b11_01_00;
        sprite_memory[380] = 6'b11_01_00;
        sprite_memory[381] = 6'b11_01_00;
        sprite_memory[382] = 6'b00_00_00;
        sprite_memory[383] = 6'b00_00_00;
        sprite_memory[384] = 6'b00_00_00;
        sprite_memory[385] = 6'b00_00_00;
        sprite_memory[386] = 6'b11_01_00;
        sprite_memory[387] = 6'b11_01_00;
        sprite_memory[388] = 6'b11_01_00;
        sprite_memory[389] = 6'b11_01_00;
        sprite_memory[390] = 6'b11_01_00;
        sprite_memory[391] = 6'b11_01_00;
        sprite_memory[392] = 6'b11_01_00;
        sprite_memory[393] = 6'b11_01_00;
        sprite_memory[394] = 6'b11_01_00;
        sprite_memory[395] = 6'b11_01_00;
        sprite_memory[396] = 6'b00_00_00;
        sprite_memory[397] = 6'b11_01_00;
        sprite_memory[398] = 6'b11_01_00;
        sprite_memory[399] = 6'b11_01_00;
        sprite_memory[400] = 6'b11_01_00;
        sprite_memory[401] = 6'b11_01_00;
        sprite_memory[402] = 6'b11_01_00;
        sprite_memory[403] = 6'b11_01_00;
        sprite_memory[404] = 6'b11_01_00;
        sprite_memory[405] = 6'b11_01_00;
        sprite_memory[406] = 6'b11_01_00;
        sprite_memory[407] = 6'b11_01_00;
        sprite_memory[408] = 6'b11_01_00;
        sprite_memory[409] = 6'b11_01_00;
        sprite_memory[410] = 6'b11_01_00;
        sprite_memory[411] = 6'b11_01_00;
        sprite_memory[412] = 6'b11_01_00;
        sprite_memory[413] = 6'b00_00_00;
        sprite_memory[414] = 6'b00_00_00;
        sprite_memory[415] = 6'b00_00_00;
        sprite_memory[416] = 6'b00_00_00;
        sprite_memory[417] = 6'b00_00_00;
        sprite_memory[418] = 6'b11_01_00;
        sprite_memory[419] = 6'b11_01_00;
        sprite_memory[420] = 6'b11_01_00;
        sprite_memory[421] = 6'b11_01_00;
        sprite_memory[422] = 6'b11_01_00;
        sprite_memory[423] = 6'b11_01_00;
        sprite_memory[424] = 6'b11_01_00;
        sprite_memory[425] = 6'b11_01_00;
        sprite_memory[426] = 6'b11_01_00;
        sprite_memory[427] = 6'b11_01_00;
        sprite_memory[428] = 6'b11_01_00;
        sprite_memory[429] = 6'b11_01_00;
        sprite_memory[430] = 6'b11_01_00;
        sprite_memory[431] = 6'b11_01_00;
        sprite_memory[432] = 6'b11_01_00;
        sprite_memory[433] = 6'b11_01_00;
        sprite_memory[434] = 6'b11_01_00;
        sprite_memory[435] = 6'b11_01_00;
        sprite_memory[436] = 6'b11_01_00;
        sprite_memory[437] = 6'b11_01_00;
        sprite_memory[438] = 6'b11_01_00;
        sprite_memory[439] = 6'b11_01_00;
        sprite_memory[440] = 6'b11_01_00;
        sprite_memory[441] = 6'b11_01_00;
        sprite_memory[442] = 6'b11_01_00;
        sprite_memory[443] = 6'b11_01_00;
        sprite_memory[444] = 6'b11_01_00;
        sprite_memory[445] = 6'b11_01_00;
        sprite_memory[446] = 6'b00_00_00;
        sprite_memory[447] = 6'b00_00_00;
        sprite_memory[448] = 6'b00_00_00;
        sprite_memory[449] = 6'b00_00_00;
        sprite_memory[450] = 6'b11_01_00;
        sprite_memory[451] = 6'b11_01_00;
        sprite_memory[452] = 6'b11_01_00;
        sprite_memory[453] = 6'b00_00_00;
        sprite_memory[454] = 6'b11_01_00;
        sprite_memory[455] = 6'b11_01_00;
        sprite_memory[456] = 6'b11_01_00;
        sprite_memory[457] = 6'b11_01_00;
        sprite_memory[458] = 6'b00_00_00;
        sprite_memory[459] = 6'b11_01_00;
        sprite_memory[460] = 6'b11_01_00;
        sprite_memory[461] = 6'b11_01_00;
        sprite_memory[462] = 6'b11_01_00;
        sprite_memory[463] = 6'b11_01_00;
        sprite_memory[464] = 6'b11_01_00;
        sprite_memory[465] = 6'b11_01_00;
        sprite_memory[466] = 6'b11_01_00;
        sprite_memory[467] = 6'b11_01_00;
        sprite_memory[468] = 6'b11_01_00;
        sprite_memory[469] = 6'b11_01_00;
        sprite_memory[470] = 6'b11_01_00;
        sprite_memory[471] = 6'b11_01_00;
        sprite_memory[472] = 6'b00_00_00;
        sprite_memory[473] = 6'b11_01_00;
        sprite_memory[474] = 6'b11_01_00;
        sprite_memory[475] = 6'b11_01_00;
        sprite_memory[476] = 6'b11_01_00;
        sprite_memory[477] = 6'b00_00_00;
        sprite_memory[478] = 6'b00_00_00;
        sprite_memory[479] = 6'b00_00_00;
        sprite_memory[480] = 6'b00_00_00;
        sprite_memory[481] = 6'b11_01_00;
        sprite_memory[482] = 6'b11_01_00;
        sprite_memory[483] = 6'b11_01_00;
        sprite_memory[484] = 6'b11_01_00;
        sprite_memory[485] = 6'b11_01_00;
        sprite_memory[486] = 6'b11_01_00;
        sprite_memory[487] = 6'b11_01_00;
        sprite_memory[488] = 6'b11_01_00;
        sprite_memory[489] = 6'b11_01_00;
        sprite_memory[490] = 6'b10_01_01;
        sprite_memory[491] = 6'b00_00_00;
        sprite_memory[492] = 6'b11_01_00;
        sprite_memory[493] = 6'b11_01_00;
        sprite_memory[494] = 6'b11_01_00;
        sprite_memory[495] = 6'b11_01_00;
        sprite_memory[496] = 6'b11_01_00;
        sprite_memory[497] = 6'b11_01_00;
        sprite_memory[498] = 6'b11_01_00;
        sprite_memory[499] = 6'b00_00_00;
        sprite_memory[500] = 6'b11_01_00;
        sprite_memory[501] = 6'b11_01_00;
        sprite_memory[502] = 6'b11_01_00;
        sprite_memory[503] = 6'b11_01_00;
        sprite_memory[504] = 6'b10_01_01;
        sprite_memory[505] = 6'b00_00_00;
        sprite_memory[506] = 6'b11_01_00;
        sprite_memory[507] = 6'b11_01_00;
        sprite_memory[508] = 6'b11_01_00;
        sprite_memory[509] = 6'b11_01_00;
        sprite_memory[510] = 6'b00_00_00;
        sprite_memory[511] = 6'b00_00_00;
        sprite_memory[512] = 6'b00_00_00;
        sprite_memory[513] = 6'b11_01_00;
        sprite_memory[514] = 6'b11_01_00;
        sprite_memory[515] = 6'b00_00_00;
        sprite_memory[516] = 6'b11_01_00;
        sprite_memory[517] = 6'b11_01_00;
        sprite_memory[518] = 6'b11_01_00;
        sprite_memory[519] = 6'b11_01_00;
        sprite_memory[520] = 6'b11_01_00;
        sprite_memory[521] = 6'b11_01_00;
        sprite_memory[522] = 6'b10_01_01;
        sprite_memory[523] = 6'b11_01_00;
        sprite_memory[524] = 6'b11_01_00;
        sprite_memory[525] = 6'b11_01_00;
        sprite_memory[526] = 6'b11_01_00;
        sprite_memory[527] = 6'b11_01_00;
        sprite_memory[528] = 6'b11_01_00;
        sprite_memory[529] = 6'b11_01_00;
        sprite_memory[530] = 6'b11_01_00;
        sprite_memory[531] = 6'b10_01_01;
        sprite_memory[532] = 6'b00_00_00;
        sprite_memory[533] = 6'b11_01_00;
        sprite_memory[534] = 6'b11_01_00;
        sprite_memory[535] = 6'b11_01_00;
        sprite_memory[536] = 6'b10_01_01;
        sprite_memory[537] = 6'b11_01_00;
        sprite_memory[538] = 6'b11_01_00;
        sprite_memory[539] = 6'b11_01_00;
        sprite_memory[540] = 6'b11_01_00;
        sprite_memory[541] = 6'b11_01_00;
        sprite_memory[542] = 6'b11_01_00;
        sprite_memory[543] = 6'b00_00_00;
        sprite_memory[544] = 6'b00_00_00;
        sprite_memory[545] = 6'b11_01_00;
        sprite_memory[546] = 6'b11_01_00;
        sprite_memory[547] = 6'b10_01_01;
        sprite_memory[548] = 6'b00_00_00;
        sprite_memory[549] = 6'b11_01_00;
        sprite_memory[550] = 6'b11_01_00;
        sprite_memory[551] = 6'b11_01_00;
        sprite_memory[552] = 6'b11_01_00;
        sprite_memory[553] = 6'b11_01_00;
        sprite_memory[554] = 6'b11_01_00;
        sprite_memory[555] = 6'b11_01_00;
        sprite_memory[556] = 6'b11_01_00;
        sprite_memory[557] = 6'b11_01_00;
        sprite_memory[558] = 6'b11_01_00;
        sprite_memory[559] = 6'b11_01_00;
        sprite_memory[560] = 6'b11_01_00;
        sprite_memory[561] = 6'b11_01_00;
        sprite_memory[562] = 6'b11_01_00;
        sprite_memory[563] = 6'b10_01_01;
        sprite_memory[564] = 6'b11_01_00;
        sprite_memory[565] = 6'b11_01_00;
        sprite_memory[566] = 6'b11_01_00;
        sprite_memory[567] = 6'b11_01_00;
        sprite_memory[568] = 6'b11_01_00;
        sprite_memory[569] = 6'b11_01_00;
        sprite_memory[570] = 6'b11_01_00;
        sprite_memory[571] = 6'b11_01_00;
        sprite_memory[572] = 6'b11_01_00;
        sprite_memory[573] = 6'b11_01_00;
        sprite_memory[574] = 6'b11_01_00;
        sprite_memory[575] = 6'b00_00_00;
        sprite_memory[576] = 6'b00_00_00;
        sprite_memory[577] = 6'b11_01_00;
        sprite_memory[578] = 6'b11_01_00;
        sprite_memory[579] = 6'b10_01_01;
        sprite_memory[580] = 6'b11_01_00;
        sprite_memory[581] = 6'b11_01_00;
        sprite_memory[582] = 6'b11_01_00;
        sprite_memory[583] = 6'b11_01_00;
        sprite_memory[584] = 6'b11_01_00;
        sprite_memory[585] = 6'b11_01_00;
        sprite_memory[586] = 6'b11_01_00;
        sprite_memory[587] = 6'b11_01_00;
        sprite_memory[588] = 6'b11_01_00;
        sprite_memory[589] = 6'b11_01_00;
        sprite_memory[590] = 6'b11_01_00;
        sprite_memory[591] = 6'b11_01_00;
        sprite_memory[592] = 6'b11_01_00;
        sprite_memory[593] = 6'b11_01_00;
        sprite_memory[594] = 6'b11_01_00;
        sprite_memory[595] = 6'b11_01_00;
        sprite_memory[596] = 6'b11_01_00;
        sprite_memory[597] = 6'b11_01_00;
        sprite_memory[598] = 6'b11_01_00;
        sprite_memory[599] = 6'b11_01_00;
        sprite_memory[600] = 6'b11_01_00;
        sprite_memory[601] = 6'b11_01_00;
        sprite_memory[602] = 6'b11_01_00;
        sprite_memory[603] = 6'b11_01_00;
        sprite_memory[604] = 6'b00_00_00;
        sprite_memory[605] = 6'b11_01_00;
        sprite_memory[606] = 6'b11_01_00;
        sprite_memory[607] = 6'b00_00_00;
        sprite_memory[608] = 6'b00_00_00;
        sprite_memory[609] = 6'b11_01_00;
        sprite_memory[610] = 6'b11_01_00;
        sprite_memory[611] = 6'b11_01_00;
        sprite_memory[612] = 6'b11_01_00;
        sprite_memory[613] = 6'b11_01_00;
        sprite_memory[614] = 6'b11_01_00;
        sprite_memory[615] = 6'b11_01_00;
        sprite_memory[616] = 6'b11_01_00;
        sprite_memory[617] = 6'b11_01_00;
        sprite_memory[618] = 6'b11_01_00;
        sprite_memory[619] = 6'b11_01_00;
        sprite_memory[620] = 6'b11_01_00;
        sprite_memory[621] = 6'b00_00_00;
        sprite_memory[622] = 6'b11_01_00;
        sprite_memory[623] = 6'b11_01_00;
        sprite_memory[624] = 6'b11_01_00;
        sprite_memory[625] = 6'b11_01_00;
        sprite_memory[626] = 6'b11_01_00;
        sprite_memory[627] = 6'b11_01_00;
        sprite_memory[628] = 6'b11_01_00;
        sprite_memory[629] = 6'b11_01_00;
        sprite_memory[630] = 6'b11_01_00;
        sprite_memory[631] = 6'b11_01_00;
        sprite_memory[632] = 6'b11_01_00;
        sprite_memory[633] = 6'b11_01_00;
        sprite_memory[634] = 6'b11_01_00;
        sprite_memory[635] = 6'b11_01_00;
        sprite_memory[636] = 6'b11_01_00;
        sprite_memory[637] = 6'b11_01_00;
        sprite_memory[638] = 6'b11_01_00;
        sprite_memory[639] = 6'b00_00_00;
        sprite_memory[640] = 6'b00_00_00;
        sprite_memory[641] = 6'b11_01_00;
        sprite_memory[642] = 6'b11_01_00;
        sprite_memory[643] = 6'b11_01_00;
        sprite_memory[644] = 6'b11_01_00;
        sprite_memory[645] = 6'b11_01_00;
        sprite_memory[646] = 6'b11_01_00;
        sprite_memory[647] = 6'b11_01_00;
        sprite_memory[648] = 6'b11_01_00;
        sprite_memory[649] = 6'b11_01_00;
        sprite_memory[650] = 6'b11_01_00;
        sprite_memory[651] = 6'b11_01_00;
        sprite_memory[652] = 6'b11_01_00;
        sprite_memory[653] = 6'b11_01_00;
        sprite_memory[654] = 6'b11_01_00;
        sprite_memory[655] = 6'b11_01_00;
        sprite_memory[656] = 6'b11_01_00;
        sprite_memory[657] = 6'b11_01_00;
        sprite_memory[658] = 6'b11_01_00;
        sprite_memory[659] = 6'b11_01_00;
        sprite_memory[660] = 6'b11_01_00;
        sprite_memory[661] = 6'b11_01_00;
        sprite_memory[662] = 6'b11_01_00;
        sprite_memory[663] = 6'b11_01_00;
        sprite_memory[664] = 6'b11_01_00;
        sprite_memory[665] = 6'b11_01_00;
        sprite_memory[666] = 6'b00_00_00;
        sprite_memory[667] = 6'b11_01_00;
        sprite_memory[668] = 6'b11_01_00;
        sprite_memory[669] = 6'b11_01_00;
        sprite_memory[670] = 6'b11_01_00;
        sprite_memory[671] = 6'b00_00_00;
        sprite_memory[672] = 6'b00_00_00;
        sprite_memory[673] = 6'b11_01_00;
        sprite_memory[674] = 6'b11_01_00;
        sprite_memory[675] = 6'b11_01_00;
        sprite_memory[676] = 6'b11_01_00;
        sprite_memory[677] = 6'b11_01_00;
        sprite_memory[678] = 6'b11_01_00;
        sprite_memory[679] = 6'b11_01_00;
        sprite_memory[680] = 6'b11_01_00;
        sprite_memory[681] = 6'b11_01_00;
        sprite_memory[682] = 6'b11_01_00;
        sprite_memory[683] = 6'b11_01_00;
        sprite_memory[684] = 6'b11_01_00;
        sprite_memory[685] = 6'b11_01_00;
        sprite_memory[686] = 6'b11_01_00;
        sprite_memory[687] = 6'b11_01_00;
        sprite_memory[688] = 6'b11_01_00;
        sprite_memory[689] = 6'b11_01_00;
        sprite_memory[690] = 6'b11_01_00;
        sprite_memory[691] = 6'b11_01_00;
        sprite_memory[692] = 6'b11_01_00;
        sprite_memory[693] = 6'b11_01_00;
        sprite_memory[694] = 6'b11_01_00;
        sprite_memory[695] = 6'b11_01_00;
        sprite_memory[696] = 6'b11_01_00;
        sprite_memory[697] = 6'b11_01_00;
        sprite_memory[698] = 6'b10_01_01;
        sprite_memory[699] = 6'b00_00_00;
        sprite_memory[700] = 6'b11_01_00;
        sprite_memory[701] = 6'b11_01_00;
        sprite_memory[702] = 6'b11_01_00;
        sprite_memory[703] = 6'b00_00_00;
        sprite_memory[704] = 6'b00_00_00;
        sprite_memory[705] = 6'b00_00_00;
        sprite_memory[706] = 6'b11_01_00;
        sprite_memory[707] = 6'b11_01_00;
        sprite_memory[708] = 6'b11_01_00;
        sprite_memory[709] = 6'b11_01_00;
        sprite_memory[710] = 6'b11_01_00;
        sprite_memory[711] = 6'b00_00_00;
        sprite_memory[712] = 6'b11_01_00;
        sprite_memory[713] = 6'b11_01_00;
        sprite_memory[714] = 6'b11_01_00;
        sprite_memory[715] = 6'b11_01_00;
        sprite_memory[716] = 6'b11_01_00;
        sprite_memory[717] = 6'b11_01_00;
        sprite_memory[718] = 6'b11_01_00;
        sprite_memory[719] = 6'b11_01_00;
        sprite_memory[720] = 6'b00_00_00;
        sprite_memory[721] = 6'b11_01_00;
        sprite_memory[722] = 6'b11_01_00;
        sprite_memory[723] = 6'b11_01_00;
        sprite_memory[724] = 6'b00_00_00;
        sprite_memory[725] = 6'b11_01_00;
        sprite_memory[726] = 6'b11_01_00;
        sprite_memory[727] = 6'b11_01_00;
        sprite_memory[728] = 6'b11_01_00;
        sprite_memory[729] = 6'b11_01_00;
        sprite_memory[730] = 6'b10_01_01;
        sprite_memory[731] = 6'b11_01_00;
        sprite_memory[732] = 6'b11_01_00;
        sprite_memory[733] = 6'b11_01_00;
        sprite_memory[734] = 6'b00_00_00;
        sprite_memory[735] = 6'b00_00_00;
        sprite_memory[736] = 6'b00_00_00;
        sprite_memory[737] = 6'b00_00_00;
        sprite_memory[738] = 6'b11_01_00;
        sprite_memory[739] = 6'b11_01_00;
        sprite_memory[740] = 6'b11_01_00;
        sprite_memory[741] = 6'b11_01_00;
        sprite_memory[742] = 6'b11_01_00;
        sprite_memory[743] = 6'b11_01_00;
        sprite_memory[744] = 6'b11_01_00;
        sprite_memory[745] = 6'b11_01_00;
        sprite_memory[746] = 6'b11_01_00;
        sprite_memory[747] = 6'b11_01_00;
        sprite_memory[748] = 6'b11_01_00;
        sprite_memory[749] = 6'b11_01_00;
        sprite_memory[750] = 6'b11_01_00;
        sprite_memory[751] = 6'b11_01_00;
        sprite_memory[752] = 6'b10_01_01;
        sprite_memory[753] = 6'b00_00_00;
        sprite_memory[754] = 6'b11_01_00;
        sprite_memory[755] = 6'b11_01_00;
        sprite_memory[756] = 6'b11_01_00;
        sprite_memory[757] = 6'b11_01_00;
        sprite_memory[758] = 6'b11_01_00;
        sprite_memory[759] = 6'b11_01_00;
        sprite_memory[760] = 6'b11_01_00;
        sprite_memory[761] = 6'b11_01_00;
        sprite_memory[762] = 6'b11_01_00;
        sprite_memory[763] = 6'b11_01_00;
        sprite_memory[764] = 6'b11_01_00;
        sprite_memory[765] = 6'b11_01_00;
        sprite_memory[766] = 6'b00_00_00;
        sprite_memory[767] = 6'b00_00_00;
        sprite_memory[768] = 6'b00_00_00;
        sprite_memory[769] = 6'b00_00_00;
        sprite_memory[770] = 6'b00_00_00;
        sprite_memory[771] = 6'b11_01_00;
        sprite_memory[772] = 6'b11_01_00;
        sprite_memory[773] = 6'b00_00_00;
        sprite_memory[774] = 6'b11_01_00;
        sprite_memory[775] = 6'b11_01_00;
        sprite_memory[776] = 6'b11_01_00;
        sprite_memory[777] = 6'b11_01_00;
        sprite_memory[778] = 6'b11_01_00;
        sprite_memory[779] = 6'b11_01_00;
        sprite_memory[780] = 6'b11_01_00;
        sprite_memory[781] = 6'b00_00_00;
        sprite_memory[782] = 6'b11_01_00;
        sprite_memory[783] = 6'b11_01_00;
        sprite_memory[784] = 6'b10_01_01;
        sprite_memory[785] = 6'b11_01_00;
        sprite_memory[786] = 6'b11_01_00;
        sprite_memory[787] = 6'b11_01_00;
        sprite_memory[788] = 6'b11_01_00;
        sprite_memory[789] = 6'b11_01_00;
        sprite_memory[790] = 6'b11_01_00;
        sprite_memory[791] = 6'b11_01_00;
        sprite_memory[792] = 6'b11_01_00;
        sprite_memory[793] = 6'b11_01_00;
        sprite_memory[794] = 6'b11_01_00;
        sprite_memory[795] = 6'b11_01_00;
        sprite_memory[796] = 6'b11_01_00;
        sprite_memory[797] = 6'b11_01_00;
        sprite_memory[798] = 6'b11_01_00;
        sprite_memory[799] = 6'b00_00_00;
        sprite_memory[800] = 6'b00_00_00;
        sprite_memory[801] = 6'b00_00_00;
        sprite_memory[802] = 6'b00_00_00;
        sprite_memory[803] = 6'b11_01_00;
        sprite_memory[804] = 6'b11_01_00;
        sprite_memory[805] = 6'b10_01_01;
        sprite_memory[806] = 6'b00_00_00;
        sprite_memory[807] = 6'b11_01_00;
        sprite_memory[808] = 6'b11_01_00;
        sprite_memory[809] = 6'b11_01_00;
        sprite_memory[810] = 6'b11_01_00;
        sprite_memory[811] = 6'b11_01_00;
        sprite_memory[812] = 6'b11_01_00;
        sprite_memory[813] = 6'b11_01_00;
        sprite_memory[814] = 6'b11_01_00;
        sprite_memory[815] = 6'b11_01_00;
        sprite_memory[816] = 6'b11_01_00;
        sprite_memory[817] = 6'b11_01_00;
        sprite_memory[818] = 6'b11_01_00;
        sprite_memory[819] = 6'b11_01_00;
        sprite_memory[820] = 6'b11_01_00;
        sprite_memory[821] = 6'b11_01_00;
        sprite_memory[822] = 6'b00_00_00;
        sprite_memory[823] = 6'b11_01_00;
        sprite_memory[824] = 6'b11_01_00;
        sprite_memory[825] = 6'b11_01_00;
        sprite_memory[826] = 6'b11_01_00;
        sprite_memory[827] = 6'b11_01_00;
        sprite_memory[828] = 6'b11_01_00;
        sprite_memory[829] = 6'b11_01_00;
        sprite_memory[830] = 6'b11_01_00;
        sprite_memory[831] = 6'b00_00_00;
        sprite_memory[832] = 6'b00_00_00;
        sprite_memory[833] = 6'b00_00_00;
        sprite_memory[834] = 6'b00_00_00;
        sprite_memory[835] = 6'b11_01_00;
        sprite_memory[836] = 6'b11_01_00;
        sprite_memory[837] = 6'b10_01_01;
        sprite_memory[838] = 6'b11_01_00;
        sprite_memory[839] = 6'b11_01_00;
        sprite_memory[840] = 6'b11_01_00;
        sprite_memory[841] = 6'b11_01_00;
        sprite_memory[842] = 6'b11_01_00;
        sprite_memory[843] = 6'b00_00_00;
        sprite_memory[844] = 6'b11_01_00;
        sprite_memory[845] = 6'b11_01_00;
        sprite_memory[846] = 6'b11_01_00;
        sprite_memory[847] = 6'b11_01_00;
        sprite_memory[848] = 6'b11_01_00;
        sprite_memory[849] = 6'b11_01_00;
        sprite_memory[850] = 6'b11_01_00;
        sprite_memory[851] = 6'b11_01_00;
        sprite_memory[852] = 6'b11_01_00;
        sprite_memory[853] = 6'b11_01_00;
        sprite_memory[854] = 6'b10_01_01;
        sprite_memory[855] = 6'b00_00_00;
        sprite_memory[856] = 6'b11_01_00;
        sprite_memory[857] = 6'b11_01_00;
        sprite_memory[858] = 6'b11_01_00;
        sprite_memory[859] = 6'b11_01_00;
        sprite_memory[860] = 6'b11_01_00;
        sprite_memory[861] = 6'b11_01_00;
        sprite_memory[862] = 6'b11_01_00;
        sprite_memory[863] = 6'b00_00_00;
        sprite_memory[864] = 6'b00_00_00;
        sprite_memory[865] = 6'b00_00_00;
        sprite_memory[866] = 6'b11_01_00;
        sprite_memory[867] = 6'b11_01_00;
        sprite_memory[868] = 6'b11_01_00;
        sprite_memory[869] = 6'b11_01_00;
        sprite_memory[870] = 6'b11_01_00;
        sprite_memory[871] = 6'b11_01_00;
        sprite_memory[872] = 6'b11_01_00;
        sprite_memory[873] = 6'b11_01_00;
        sprite_memory[874] = 6'b11_01_00;
        sprite_memory[875] = 6'b10_01_01;
        sprite_memory[876] = 6'b00_00_00;
        sprite_memory[877] = 6'b11_01_00;
        sprite_memory[878] = 6'b11_01_00;
        sprite_memory[879] = 6'b11_01_00;
        sprite_memory[880] = 6'b11_01_00;
        sprite_memory[881] = 6'b11_01_00;
        sprite_memory[882] = 6'b11_01_00;
        sprite_memory[883] = 6'b11_01_00;
        sprite_memory[884] = 6'b11_01_00;
        sprite_memory[885] = 6'b11_01_00;
        sprite_memory[886] = 6'b10_01_01;
        sprite_memory[887] = 6'b11_01_00;
        sprite_memory[888] = 6'b11_01_00;
        sprite_memory[889] = 6'b11_01_00;
        sprite_memory[890] = 6'b11_01_00;
        sprite_memory[891] = 6'b11_01_00;
        sprite_memory[892] = 6'b00_00_00;
        sprite_memory[893] = 6'b11_01_00;
        sprite_memory[894] = 6'b11_01_00;
        sprite_memory[895] = 6'b00_00_00;
        sprite_memory[896] = 6'b00_00_00;
        sprite_memory[897] = 6'b00_00_00;
        sprite_memory[898] = 6'b00_00_00;
        sprite_memory[899] = 6'b11_01_00;
        sprite_memory[900] = 6'b11_01_00;
        sprite_memory[901] = 6'b11_01_00;
        sprite_memory[902] = 6'b11_01_00;
        sprite_memory[903] = 6'b11_01_00;
        sprite_memory[904] = 6'b11_01_00;
        sprite_memory[905] = 6'b11_01_00;
        sprite_memory[906] = 6'b11_01_00;
        sprite_memory[907] = 6'b10_01_01;
        sprite_memory[908] = 6'b11_01_00;
        sprite_memory[909] = 6'b11_01_00;
        sprite_memory[910] = 6'b11_01_00;
        sprite_memory[911] = 6'b11_01_00;
        sprite_memory[912] = 6'b11_01_00;
        sprite_memory[913] = 6'b00_00_00;
        sprite_memory[914] = 6'b11_01_00;
        sprite_memory[915] = 6'b11_01_00;
        sprite_memory[916] = 6'b11_01_00;
        sprite_memory[917] = 6'b11_01_00;
        sprite_memory[918] = 6'b11_01_00;
        sprite_memory[919] = 6'b11_01_00;
        sprite_memory[920] = 6'b11_01_00;
        sprite_memory[921] = 6'b11_01_00;
        sprite_memory[922] = 6'b11_01_00;
        sprite_memory[923] = 6'b11_01_00;
        sprite_memory[924] = 6'b10_01_01;
        sprite_memory[925] = 6'b00_00_00;
        sprite_memory[926] = 6'b11_01_00;
        sprite_memory[927] = 6'b11_01_00;
        sprite_memory[928] = 6'b00_00_00;
        sprite_memory[929] = 6'b00_00_00;
        sprite_memory[930] = 6'b11_01_00;
        sprite_memory[931] = 6'b11_01_00;
        sprite_memory[932] = 6'b11_01_00;
        sprite_memory[933] = 6'b11_01_00;
        sprite_memory[934] = 6'b11_01_00;
        sprite_memory[935] = 6'b11_01_00;
        sprite_memory[936] = 6'b11_01_00;
        sprite_memory[937] = 6'b11_01_00;
        sprite_memory[938] = 6'b11_01_00;
        sprite_memory[939] = 6'b11_01_00;
        sprite_memory[940] = 6'b11_01_00;
        sprite_memory[941] = 6'b11_01_00;
        sprite_memory[942] = 6'b11_01_00;
        sprite_memory[943] = 6'b11_01_00;
        sprite_memory[944] = 6'b11_01_00;
        sprite_memory[945] = 6'b11_01_00;
        sprite_memory[946] = 6'b11_01_00;
        sprite_memory[947] = 6'b11_01_00;
        sprite_memory[948] = 6'b11_01_00;
        sprite_memory[949] = 6'b11_01_00;
        sprite_memory[950] = 6'b11_01_00;
        sprite_memory[951] = 6'b11_01_00;
        sprite_memory[952] = 6'b11_01_00;
        sprite_memory[953] = 6'b11_01_00;
        sprite_memory[954] = 6'b11_01_00;
        sprite_memory[955] = 6'b11_01_00;
        sprite_memory[956] = 6'b10_01_01;
        sprite_memory[957] = 6'b11_01_00;
        sprite_memory[958] = 6'b11_01_00;
        sprite_memory[959] = 6'b11_01_00;
        sprite_memory[960] = 6'b00_00_00;
        sprite_memory[961] = 6'b11_01_00;
        sprite_memory[962] = 6'b11_01_00;
        sprite_memory[963] = 6'b11_01_00;
        sprite_memory[964] = 6'b11_01_00;
        sprite_memory[965] = 6'b11_01_00;
        sprite_memory[966] = 6'b11_01_00;
        sprite_memory[967] = 6'b11_01_00;
        sprite_memory[968] = 6'b11_01_00;
        sprite_memory[969] = 6'b11_01_00;
        sprite_memory[970] = 6'b11_01_00;
        sprite_memory[971] = 6'b11_01_00;
        sprite_memory[972] = 6'b11_01_00;
        sprite_memory[973] = 6'b11_01_00;
        sprite_memory[974] = 6'b11_01_00;
        sprite_memory[975] = 6'b11_01_00;
        sprite_memory[976] = 6'b11_01_00;
        sprite_memory[977] = 6'b11_01_00;
        sprite_memory[978] = 6'b11_01_00;
        sprite_memory[979] = 6'b11_01_00;
        sprite_memory[980] = 6'b11_01_00;
        sprite_memory[981] = 6'b11_01_00;
        sprite_memory[982] = 6'b11_01_00;
        sprite_memory[983] = 6'b11_01_00;
        sprite_memory[984] = 6'b11_01_00;
        sprite_memory[985] = 6'b11_01_00;
        sprite_memory[986] = 6'b11_01_00;
        sprite_memory[987] = 6'b11_01_00;
        sprite_memory[988] = 6'b11_01_00;
        sprite_memory[989] = 6'b11_01_00;
        sprite_memory[990] = 6'b11_01_00;
        sprite_memory[991] = 6'b11_01_00;
        sprite_memory[992] = 6'b00_00_00;
        sprite_memory[993] = 6'b11_01_00;
        sprite_memory[994] = 6'b11_01_00;
        sprite_memory[995] = 6'b11_01_00;
        sprite_memory[996] = 6'b11_01_00;
        sprite_memory[997] = 6'b11_01_00;
        sprite_memory[998] = 6'b11_01_00;
        sprite_memory[999] = 6'b11_01_00;
        sprite_memory[1000] = 6'b11_01_00;
        sprite_memory[1001] = 6'b11_01_00;
        sprite_memory[1002] = 6'b11_01_00;
        sprite_memory[1003] = 6'b11_01_00;
        sprite_memory[1004] = 6'b11_01_00;
        sprite_memory[1005] = 6'b11_01_00;
        sprite_memory[1006] = 6'b11_01_00;
        sprite_memory[1007] = 6'b11_01_00;
        sprite_memory[1008] = 6'b11_01_00;
        sprite_memory[1009] = 6'b11_01_00;
        sprite_memory[1010] = 6'b11_01_00;
        sprite_memory[1011] = 6'b11_01_00;
        sprite_memory[1012] = 6'b11_01_00;
        sprite_memory[1013] = 6'b11_01_00;
        sprite_memory[1014] = 6'b11_01_00;
        sprite_memory[1015] = 6'b11_01_00;
        sprite_memory[1016] = 6'b11_01_00;
        sprite_memory[1017] = 6'b11_01_00;
        sprite_memory[1018] = 6'b11_01_00;
        sprite_memory[1019] = 6'b11_01_00;
        sprite_memory[1020] = 6'b11_01_00;
        sprite_memory[1021] = 6'b11_01_00;
        sprite_memory[1022] = 6'b11_01_00;
        sprite_memory[1023] = 6'b11_01_00;
    end

    always @(posedge clk) begin
        pixel_color <= sprite_memory[pixel_index]; 
    end

endmodule